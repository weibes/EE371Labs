/*
module collisionDetector (Clock, reset, normalCollisionDetected, endCollisionDetected, collisionRequest, playerPieceX,
								  playerPieceY, playerPieceOffsets, staticPiecesAddr, staticPiecesRow);
	input logic Clock, reset, collisionRequest;
	input logic [5:0] playerPiecesOffsets;
	input logic [11:0] staticPiecesRow;
	input logic [4:0] playerPieceY, playerPieceX;
	
	output logic collisionReady, normalCollisionDetected, endCollisionDetected
	
	
endmodule
*/