module displayDriver(dataIn, Clock, Reset,  VGA_R, VGA_G, VGA_B, VGA_BLANK_N, VGA_CLK, VGA_HS, VGA_SYNC_N, VGA_VS);
	input logic [39:0] dataIn [9:0];
	input logic Clock, Reset;
	
	output [7:0] VGA_R;
	output [7:0] VGA_G;
	output [7:0] VGA_B;
	output VGA_BLANK_N;
	output VGA_CLK;
	output VGA_HS;
	output VGA_SYNC_N;
	output VGA_VS;
	
	
	enum {draw_board, game_play, game_over} ps, ns;
	
	
	
	always_comb begin
		case (ps)
			draw_board:	if (
	
	end // always_comb begin
	
	
	always_ff @(posedge Clock) begin
		
	
	end // always_ff @(posedge Clock) begin
	
	
	VGA_framebuffer fb (
		.clk50			(clock), 
		.reset			(1'b0), 
		.x(finalX), 
		.y(finalY),
		.pixel_color(pixel_color && KEY[1]), 
		.pixel_write	(1'b1),
		.VGA_R, 
		.VGA_G, 
		.VGA_B, 
		.VGA_CLK, 
		.VGA_HS, 
		.VGA_VS,
		.VGA_BLANK_n	(VGA_BLANK_N), 
		.VGA_SYNC_n		(VGA_SYNC_N));
		
		
	
endmodule

